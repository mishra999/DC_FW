library IEEE;
    use IEEE.STD_LOGIC_1164.ALL;
    use IEEE.NUMERIC_STD.ALL;
    use IEEE.STD_LOGIC_MISC.ALL;
    use IEEE.STD_LOGIC_UNSIGNED.ALL;
library unisim;
    use unisim.vcomponents.all;
library unimacro;
    use unimacro.vcomponents.all;
Library work;
    use work.klm_scint_pkg.all;
    -- use work.conc_intfc_pkg.all;
    -- use work.klm_scrod_pkg.all;
    -- use work.tdc_pkg.all;

--!
--!### Operation of WaveformReadout module:
--!    <p>The job of this module is to manage all the modules needed for waveform
--!readout, pedestal management,  and feature extraction.
--!When a local trigger is received, the region of interest is calculated
--!and the trigger is put into the queue. If the queue gets too full, the next 
--!packets will be of the 'simple' type to speed things up, otherwise digitization
--!will proceed</p>
--!    <p>The FSM ro_states starts digitization and ultimately sends DAQ packets.
--!Digitization and processing happens in parallel on both busses.
--!This is taken care of by each SingleBusProcessing module. In each
--!of these modules, TrigBit2Mask modules generate one channel mask for
--!each ASIC on the bus. The module DigitizeAndShiftOutData begins
--!digitizing the first window for all ASICs on the bus, and meanwhile,
--!PedFetchQueue starts fetching pedestals for the hit channel which is first
--!to be shifted out. The ped fetcher arbitrates which bus (A/B) gets RAM
--!access first.</p>
--!    <p>As digitization of the first window finishes, all channels on any
--!hit ASICs shift out 32 samples** in parallel. ThresholdCheck writes all
--!hit channels to their own deticated FIFO in WaveAndPedStaging while at
--!the same time checking each channel to see if it crossed a programable
--!threshold value. Digitization of the remaining windows in the ROI
--!follows suit. When finished shifting out the last window, the new channel
--!mask generated by ThresholdCheck is used to flush stale jobs from the
--!PedFetchQueue and tell ProcWaveform which channels to process.</p>
--!<p>As ProcWaveform finishes its first job, it tries to send the results
--!to ro_states. An arbiter prevents collisions in case both buses
--!finish at the same time. ro_states keeps track of first hit, last
--!hit, and resets all the FIFOs when the event is finished.</p>
--!    <p>For pedestal measurement and writing, ped_sub_ena must be high,
--! then force_trig initiates the process. MeasurePeds keeps an eye
--! on the window counter and triggers readout only after it has passed.
--! in this mode, the wave and ped FIFOs in WaveAndPedStaging are taken over
--! and used to make a 24-bit wide summation. After 2**N_BITS_AVG_g dig cycles,
--! the averaged pedestals are shifted out and written to SRAM</p>
--!    <p>Lastly, two debug tools have been included in this firmeare.
--!Debug waveforms are written to a fifo every time a waveform is processessed.
--!This FIFO just fills up until somebody reads it from the register interface.
--!The second is a histogram of charge measurements done using BRAM. It fills
--!continuously until someone issues a reset</p>
--!
--!### DAQ Packet Format
--!| Word   |              Word contents                  |
--!|--------|---------------------------------------------|
--!| 1      |<pre>type(2:0) / lane(4:0) / axis(0) / chnl(6:0) </pre>|
--!| 2      |<pre>                  ctime(15:0)               </pre>|
--!| 3      |<pre>SIMP / TB5 /              TDC(13:0)         </pre>|
--!| 4      |<pre>TBD(3:0)   /              chg(11:0)         </pre>|
--!

-- #### Deficiencies:
--1. For now, we shift out whole windows only, if we calculate a finer ROI,
--then we can perhaps shift out fewer samples to save time.

entity WaveformReadout is
    generic (
        nominal_LE_sample_number_g: std_logic_vector(13 downto 0) := "00000000001000";
        FORCE_TRIG_BUF_DEPTH_g    : integer := 6;
        TRG_BUFF_DEPTH_g          : integer := 4;
        TRIG_QUEUE_DEPTH_g        : integer := 15;
        -- TQ_PROG_FULL_THRESH_g     : integer := 3;
        CALC_ROI_LAG_g            : integer := 2;
        T_WAIT_2C_IF_QUEUE_FULL_g : integer := 31; -- tried 6 and got all zeros from TARGETX, yet fine in sim -- maybe try as register
        reset_buff_depth_g        : integer := 10;
        SLC_STAT_BUFF_DEPTH_g     : integer := 4;
        packet_type_g             : std_logic_vector(7 downto 0):= X"80"; -- marks scintillators hits for DataConcentrator
        LAST_WINDOW_ADDRESS       : std_logic_vector(8 downto 0) := "111111111";
        N_BITS_AVG_g              : integer := 7;
        T_wait_busy_to_come_up_g  : integer := 31;
        -- FINE_LOOKBACK_g           : std_logic_vector(10 downto 0) := "00000000000"; -- 1 clk period resolution
        USE_PULSE_HEIGHT_HIST     : std_logic := '0';
        USE_DBG_WAVE_FIFO         : std_logic := '0';
        max_proc_time_g           : std_logic_vector(15 downto 0) := "0011000110011100" -- 100us
    );
    port (
        -- main inputs
        clk                   : in  std_logic := '0';
        busy                  : out std_logic;
        b2tt_runreset         : in  std_logic := '0';
        trig                  : in  trig_info_type_0 := null_trig_info_t0;

        -- signals with SamplingLgc
        ana_wr_ena_mask       : out TARGETX_analong_wr_ena_mask_t;
        
        -- signals with HitDataSerializer
        localtrg              : in  std_logic := '0';
        ped_meas_start        : in  std_logic := '0';
        sps_reset             : in  std_logic := '0';
        cur_win               : in  std_logic_vector(8 downto 0);
        
        -- nxt                   : in  std_logic := '0';
        -- tbfifo_rden           : out  std_logic_vector(9 downto 0);
      --! daq data ports
        qt_fifo_rd_en         : in  std_logic := '0';
        qt_fifo_dout          : out std_logic_vector (17 downto 0);
        qt_fifo_empty         : out std_logic;
        qt_fifo_err_cnt       : out std_logic_vector(15 downto 0); -- counter for daq data fifo overflows
        qt_fifo_evt_rdy       : out std_logic;
        full_proc_cnt         : out std_logic_vector(15 downto 0);
        simp_proc_cnt         : out std_logic_vector(15 downto 0);
        null_proc_cnt         : out std_logic_vector(15 downto 0);

        -- pedestal RAM access
        RAM_IO                : inout std_logic_vector(7 downto 0) := (others => '0');
        RAM_WEb               : out std_logic;
        RAM_OEb               : out std_logic;
        RAM_ADDR              : out std_logic_vector(21 downto 0);

        -- BusA signals
        BUSA_DO               : in  std_logic_vector(14 downto 0) := (others => '0');
        BUSA_RAMP             : out std_logic;
        BUSA_CLR              : out std_logic;
        BUSA_RD_COLSEL        : out std_logic_vector(5 downto 0);
        BUSA_RD_ENA           : out std_logic;
        BUSA_RD_ROWSEL        : out std_logic_vector(2 downto 0);
        BUSA_SAMPLESEL        : out std_logic_vector(4 downto 0);
        BUSA_SR_CLEAR         : out std_logic;
        BUSA_SR_SEL           : out std_logic;

        -- BusB signals
        BUSB_DO               : in  std_logic_vector(14 downto 0) := (others => '0');
        BUSB_RAMP             : out std_logic;
        BUSB_CLR              : out std_logic;
        BUSB_RD_COLSEL        : out std_logic_vector(5 downto 0);
        BUSB_RD_ENA           : out std_logic;
        BUSB_RD_ROWSEL        : out std_logic_vector(2 downto 0);
        BUSB_SAMPLESEL        : out std_logic_vector(4 downto 0);
        BUSB_SR_CLEAR         : out std_logic;
        BUSB_SR_SEL           : out std_logic;

        -- TargetX DC signals
        SAMPLESEL_ANY         : out std_logic_vector(9 downto 0);
        SR_CLOCK              : out std_logic_vector(9 downto 0);

        -- SCROD config registers
        wave_config           : in wave_config_t := default_wave_config;

        -- status registers
        wave_stat             : out waveform_stat_t := wave_stat_0;
        debug_wave_we         : out std_logic_vector(1 downto 0);
        debug_wave_din        : out slv12(1 downto 0);
        SPS_hist_rd_data      : out slv16(1 downto 0)
    );
end WaveformReadout;


architecture Behavioral of WaveformReadout is

    type trig_staging_FSM is (IDLE, WAIT_VALID, PROCESSING_REQ, WAIT_ACK);
    type modify_sampling_mask_FSM is (IDLE, WAIT_DONE);
    type ro_states is (IDLE, WAIT_RESET, CHECK_VALID, WAIT_WAVEFORM_READOUT, SEND_HITS, CHECK_DONE, STOP, SEND_SIMPLE);


--SYNCHRONOUS SIGNALS BY PROCESS WHICH DRIVES THEM
 
    --! ppln_stat: 
    signal wave_stat_i : wave_stat_vec(SLC_STAT_BUFF_DEPTH_g - 1 downto 0) := (others => wave_stat_0);

    --! conf_dffs:
    signal wave_config_q1 : wave_config_t := default_wave_config;
    signal wave_config_q2 : wave_config_t := default_wave_config;
    signal wave_config_q3 : wave_config_t := default_wave_config;
    signal wave_config_q4 : wave_config_t := default_wave_config;
    signal wave_config_q5 : wave_config_t := default_wave_config;
    signal wave_config_q6 : wave_config_t := default_wave_config;

    --! rst_buff:
    signal i_b2tt_runreset : std_logic_vector(reset_buff_depth_g - 1 downto 0);
    signal single_bus_reset_q1      : std_logic := '0';

    --! busy_lgc:
    signal or_busy_sr           : std_logic_vector(5 downto 0) := (others => '0');
    -- signal either_bus_busy     : std_logic := '0';

    --! trg_buff:
    signal i_localtrg : std_logic_vector(TRG_BUFF_DEPTH_g - 1 downto 0);

    --! ped_meas_start_buffer:
    signal ped_meas_start_sr : std_logic_vector(FORCE_TRIG_BUF_DEPTH_g-1 downto 0) := (others => '0');
    signal sps_reset_sr  : std_logic_vector(FORCE_TRIG_BUF_DEPTH_g-1 downto 0) := (others => '0');

    --! SRAM_mux:
    signal meas_peds_ena       : std_logic;
    signal i_N_readout_samples : std_logic_vector(8 downto 0) := "000011111";
    signal i_RAM_WEb           : std_logic := '1';
    signal i_RAM_din           : std_logic_vector(7 downto 0) := (others => '0');
    signal RAM_din             : std_logic_vector(7 downto 0) := (others => '0');
    signal RAM_rw              : std_logic := '1';

    --! ena_logic:
    signal single_bus_ena    : std_logic := '0';
    signal SPS_measure_start : std_logic_vector(1 downto 0) := "00";

    --! asic_chan_win_mux:
    signal i_trig_bits       : slv5(9 downto 0) := (others=>(others=>'0'));
    signal starting_win_samp : slv14(9 downto 0) := (others => (others=>'0'));
    signal LE_ctime          : slv14(9 downto 0) := (others => (others=>'0'));
    signal first_dig_win     : std_logic_vector(8 downto 0) := (others=>'0');
    signal last_dig_win      : std_logic_vector(8 downto 0) := (others=>'0');
    signal asic_mask         : std_logic_vector(9 downto 0) := (others => '0');

    --! trg_proc:
    signal trig_staging      : trig_staging_FSM := IDLE;
    signal trig_in_t0        : trig_info_type_0 := null_trig_info_t0; --! copy of input trig without ROI
    signal trg_stg_fsm_ctr   : integer range 0 to (CALC_ROI_LAG_g + N_ASICS) := 0;
    signal calc_roi_ena      : std_logic := '0';
    signal trg_proc_busy     : std_logic := '0';
    signal mask_windows      : std_logic := '0';
    signal trig_queue_wr_ena : std_logic := '0';

    --! trg_queue:
    signal wr_ptr             : integer range 0 to TRIG_QUEUE_DEPTH_g - 1 := 0;
    signal rd_ptr             : integer range 0 to TRIG_QUEUE_DEPTH_g - 1 := 0;
    signal wr_ptr_nxt         : integer range 0 to TRIG_QUEUE_DEPTH_g - 1 := 0;
    signal rd_ptr_nxt         : integer range 0 to TRIG_QUEUE_DEPTH_g - 1 := 0;
    signal queue_empty        : std_logic := '1';
    -- signal queue_above_thresh : std_logic := '0';
    -- signal queue_getting_full : std_logic := '0';
    signal queue_full         : std_logic := '0';
    signal start_readout      : std_logic := '0';
    signal trig_queue         : trig_queue_type(TRIG_QUEUE_DEPTH_g - 1 downto 0) := (others => null_trig_info_t1); -- triggers on deck
    signal trig_q0            : trig_info_type_1 := null_trig_info_t1;                               

    --! mask_unmask_proc:
    signal modify_sampling_mask  : modify_sampling_mask_FSM := IDLE;
    signal mod_samp_msk_fsm_ctr  : integer range 0 to 3 := 0;
    signal mask_ack              : std_logic := '0';
    signal unmask_ack            : std_logic := '0';
    signal i_ana_wr_ena_mask     : TARGETX_analong_wr_ena_mask_t := null_TX_ana_wr_ena_mask;
    
    --! hit_bldr:
    signal ro_state             : ro_states := IDLE;
    signal ro_st_fsm_ctr        : integer range 0 to T_WAIT_2C_IF_QUEUE_FULL_g := 0;
    signal i_last_hit           : std_logic_vector(1 downto 0) := "00";
    signal i_first_hit          : std_logic := '1';
    signal simple_mode_ena      : std_logic := '0';
    signal proc_queue_quick     : std_logic := '0';
    signal hit_bldr_fsm_busy    : std_logic := '0';
    signal ro_reset             : std_logic := '0';
    signal daq_axis_i           : std_logic := '0';
    signal daq_chan_i           : std_logic_vector(6 downto 0) := (others => '0');
    signal daq_chan_base        : std_logic_vector(6 downto 0) := (others => '0');
    signal trig_bits_i          : std_logic_vector(4 downto 0) := (others => '0');
    signal simp                 : std_logic := '0';
    -- signal le_time_c            : std_logic_vector(8 downto 0) := (others => '0');
    -- signal le_time_f            : std_logic_vector(4 downto 0) := (others => '0');
    signal le_time_i            : std_logic_vector(13 downto 0) := (others => '0');
    signal L0_ctime_i           : std_logic_vector(15 downto 0) := (others => '0');
    signal peak_i               : std_logic_vector(11 downto 0) := (others => '0');
    signal daq_start_ro         : std_logic := '0';
    signal i_full_proc_cnt      : std_logic_vector(15 downto 0) := (others => '0');
    signal i_simp_proc_cnt      : std_logic_vector(15 downto 0) := (others => '0');
    signal i_null_proc_cnt      : std_logic_vector(15 downto 0) := (others => '0');
    signal daq_asic_mask        : std_logic_vector(9 downto 0) := (others => '0');
    signal simp_asic_mask       : std_logic_vector(9 downto 0) := (others => '0');
    signal unmask_windows       : std_logic := '0';
    signal rx_features_ack      : std_logic_vector(1 downto 0) := (others => '0');
    signal ser_run_q0           : std_logic := '0';
    signal HitData_i            : KlmScrodHitDataType := KlmScrodHitDataNull;
   
    --! ppln_hit_data:
    signal ser_run_q1           : std_logic := '0';
    signal ser_run_q2           : std_logic := '0';
    signal ser_run_q3           : std_logic := '0';
    signal HitData  : KlmScrodHitDataType := KlmScrodHitDataNull;

 

--! ASYNCHRONOUSLY DRIVEN SIGNALS
    signal single_bus_reset  : std_logic := '0';
    signal disambig_tb5      : std_logic := '1';
    -- signal or_busy_status    : std_logic := '0';
    -- signal L0_ctime_win      : slv11(9 downto 0) := (others=>(others=>'0'));

-- SIGNALS DRIVEN BY INSTANTIATED ENTITIES

    --! CALC_ROI:
    signal trig_in_t1    : trig_info_type_1 := null_trig_info_t1; -- copy of input trig with ROI added


    --! busA/busB:
    signal i_ped_fetch_asic_no : slv3(1 downto 0);-- := (others => "000");
    signal ped_fetch_chan      : slv4(1 downto 0) := (others => "0000");
    signal ped_win_samp_start  : slv14(1 downto 0) := (others=>(others=>'0'));
    signal ped_fetch_ena       : std_logic_vector(1 downto 0) := (others => '0');
    signal BUSA_WINSEL         : std_logic_vector(8 downto 0) := (others => '0');
    signal BUSB_WINSEL         : std_logic_vector(8 downto 0) := (others => '0');
    signal rx_features_ena     : std_logic_vector(1 downto 0) := (others => '0');
    signal last_hit            : std_logic_vector(1 downto 0) := "00";
    signal peak              : slv12(1 downto 0) := (others => "000000000000");
    signal le_time             : slv9(1 downto 0) := (others => "000000000");
    signal daq_chan            : slv7(1 downto 0) := (others => "0000000");
    signal daq_asic            : i5(1 downto 0) := (0, 0);
    -- signal DigStoreProcBusy    : std_logic_vector(1 downto 0) := "00";
    signal DigNShiftBusy       : std_logic_vector(1 downto 0) := "00";
    -- signal DigBusy             : std_logic_vector(1 downto 0) := "00";
    signal ShiftOutWinBusy     : std_logic_vector(1 downto 0) := "00";
    signal ShiftOutSampBusy    : std_logic_vector(1 downto 0) := "00";
    -- signal FeatExtBusy         : std_logic_vector(1 downto 0) := "00";
    -- signal PedFetchQueueBusy   : std_logic_vector(1 downto 0) := "00";
    signal avg_peds_busy       : std_logic_vector(1 downto 0) := "00";
    signal wr_peds2sram_ena    : std_logic_vector(1 downto 0) := (others=>'0');
    signal even_sample         : slv12(1 downto 0) := (others => (others=>'0'));
    signal odd_sample          : slv12(1 downto 0) := (others => (others=>'0'));
    signal sram_asic_addr      : slv3(1 downto 0) := (others=>(others=>'0'));
    signal sram_chan_addr      : slv4(1 downto 0) := (others=>(others=>'0'));
    signal sram_samp_addr      : slv4(1 downto 0) := (others=>(others=>'0'));

    --! ped_fetcher:
    signal ped_fetch_ack       : std_logic_vector(1 downto 0) := (others => '0');
    signal ped_fifo_asic_sel   : std_logic_vector(4 downto 0) := (others => '0');
    signal ped_fifo_chan_sel   : std_logic_vector(3 downto 0) := (others => '0');
    signal ped_fifo_wr_ena     : std_logic_vector(1 downto 0) := (others => '0');
    signal ped_fifo_din        : std_logic_vector(11 downto 0) := (others => '0');
    signal RAM_rd_addr         : std_logic_vector(21 downto 0) := (others => '1');

    --! ped_writer:
    signal RAM_wr_addr      : std_logic_vector(21 downto 0) := (others => '1');
    signal wr_peds2sram_ack : std_logic_vector(1 downto 0) := (others=>'0');

    --! ped_measure:
    signal ped_meas_win         : std_logic_vector(8 downto 0) := (others=>'0');
    signal ped_start_ro         : std_logic := '0';
    signal prime_fifos          : std_logic := '0';
    signal avg_peds_ena         : std_logic := '0';
    signal summing_ena          : std_logic := '0';

    -- HitData_Serializer_i :
    signal ser_busy     : std_logic := '0';
    
    --! sda_buff:
    signal RAM_do :  std_logic_vector(7 downto 0) := (others => '0');

begin

------------------- ASYNCHRONOUS LOGIC ---------------------------------------------

    single_bus_reset <= ro_reset; -- or rst_from_sps_fsm;
    BUSA_RD_ROWSEL <= BUSA_WINSEL(2 downto 0); -- Kurtis says bit pattern is more complicated...
    BUSB_RD_ROWSEL <= BUSB_WINSEL(2 downto 0); -- ...may be shuffled in UCF or elsewhere in firmware
    -- BUSA_RD_ROWSEL <= BUSA_WINSEL(1) & BUSA_WINSEL(2) & BUSA_WINSEL(0);
    -- BUSB_RD_ROWSEL <= BUSB_WINSEL(1) & BUSB_WINSEL(2) & BUSB_WINSEL(0);
    BUSA_RD_COLSEL <= BUSA_WINSEL(8 downto 3);
    BUSB_RD_COLSEL <= BUSB_WINSEL(8 downto 3);
    -- dbg_start_ro <= (force_trig_sr(force_trig_sr'left) and not (wave_config_q6.measure_peds or wave_config_q6.use_loop_trig));
    -- asic_chan_win_sel <= wave_config_q6.measure_peds & wave_config_q6.use_ftsw_trig;
    -- bus_mask <= daq_bus_mask or ped_bus_mask;
    ana_wr_ena_mask <= i_ana_wr_ena_mask;
    trig_in_t1.L0_ctime <= trig_in_t0.L0_ctime;
    trig_in_t1.ana_addr <= trig_in_t0.ana_addr;
    trig_in_t1.mask <= trig_in_t0.mask;
    trig_in_t1.L1_ctime <= trig_in_t0.L1_ctime;
    trig_in_t1.bits <= trig_in_t0.bits;
    wave_stat_i(0).fe_dbg_a <= ShiftOutSampBusy(0) & ShiftOutWinBusy(0);
    wave_stat_i(0).fe_dbg_b <= ShiftOutSampBusy(1) & ShiftOutWinBusy(1);
    -- or_busy_status <= or_reduce(DigStoreProcBusy)
    --                   or or_reduce(DigNShiftBusy)
    --                   or or_reduce(DigBusy)
    --                   or or_reduce(ShiftOutWinBusy)
    --                   or or_reduce(ShiftOutSampBusy)
    --                   or or_reduce(FeatExtBusy)
    --                   or or_reduce(PedFetchQueueBusy);
    -- trg_proc_cnt <= i_trg_proc_cnt(31 downto 24) & i_trg_proc_cnt(7 downto 0); 
    full_proc_cnt <= i_full_proc_cnt;
    simp_proc_cnt <= i_simp_proc_cnt;
    null_proc_cnt <= i_null_proc_cnt;
    -- or_calc_roi_busy <= or_reduce(calc_roi_busy);
    disambig_tb5 <= wave_config_q6.use_ftsw_trig;
    -- gen_calcROI_windows : for i in 0 to 9 generate
    --     L0_ctime_win(i) <= trig_in_t0.L0_ctime(i)(10 downto 0);
    -- end generate;
        
--------------------- SYNCHRONOUS LOGIC ---------------------------------------------

    ppln_stat: process(clk, wave_stat_i)
    begin
        wave_stat <= wave_stat_i(wave_stat_i'left);
        wave_stat_i(wave_stat_i'left downto 1) <= wave_stat_i(wave_stat_i'left - 1 downto 0);
    end process;
    
    conf_dffs: process(clk, wave_config, wave_config_q1, wave_config_q2,
                       wave_config_q3, wave_config_q4, wave_config_q5)
    begin
        if rising_edge(clk) then
            wave_config_q1 <= wave_config;
            wave_config_q2 <= wave_config_q1;
            wave_config_q3 <= wave_config_q2;
            wave_config_q4 <= wave_config_q3;
            wave_config_q5 <= wave_config_q4;
            wave_config_q6 <= wave_config_q5;
        end if;
    end process conf_dffs;

    rst_buff: process(clk, b2tt_runreset, i_b2tt_runreset)
    begin
        if rising_edge(clk) then
            i_b2tt_runreset(reset_buff_depth_g - 1 downto 1) <= i_b2tt_runreset(reset_buff_depth_g - 2 downto 0);
            i_b2tt_runreset(0) <= b2tt_runreset;
            single_bus_reset_q1 <= single_bus_reset;
        end if;
    end process rst_buff;


    busy_lgc: process(clk, DigNShiftBusy, queue_full)
    begin
        if rising_edge(clk) then
            -- or_busy_sr <= or_busy_sr(or_busy_sr'left - 1 downto 0) & or_busy_status;
            or_busy_sr <= or_busy_sr(or_busy_sr'left - 1 downto 0) & or_reduce(DigNShiftBusy);
            -- either_bus_busy <= or_busy_sr(or_busy_sr'left);
            wave_stat_i(0).wave_proc_busy <= hit_bldr_fsm_busy;
            -- busy <= localtrg or calc_roi_busy(0) or calc_roi_busy(1) or queue_full;
            busy <= trg_proc_busy or queue_full;
        end if;
    end process busy_lgc;
    
    
    trg_buff: process(clk, localtrg)
    begin
        if rising_edge(clk) then
            i_localtrg <= i_localtrg(i_localtrg'left - 1 downto 0) & localtrg;
        end if;
    end process;
    

    ped_meas_start_buffer: process(clk, ped_meas_start)
    begin
        if rising_edge(clk) then
            ped_meas_start_sr <= ped_meas_start_sr(ped_meas_start_sr'left - 1 downto 0) & ped_meas_start;
        end if;
    end process;
    
    
    sps_reset_buffer: process(clk, sps_reset)
    begin
        if rising_edge(clk) then
            sps_reset_sr <= sps_reset_sr(sps_reset_sr'left - 1 downto 0) & sps_reset;
        end if;
    end process;
    
    
    ----------------------------------------------------------------------------
    -- ADDRESS MULTIPLEXER AND PIPELINE FOR SRAM CONTROL --
    ----------------------------------------------------------------------------
    SRAM_mux: process (clk, wave_config_q6.measure_peds, ped_meas_start_sr, i_RAM_din,
            RAM_wr_addr, RAM_rd_addr, i_RAM_WEb)
    begin
        if rising_edge(clk) then
            RAM_din  <= i_RAM_din; -- DFF for matching phase with address
            RAM_WEb <= i_RAM_WEb; -- DFF for matching phase with address
            if wave_config_q6.measure_peds = '1' then
                RAM_rw <= '0';
                RAM_OEb <= '1';
                RAM_ADDR <= RAM_wr_addr;
                meas_peds_ena <= ped_meas_start_sr(ped_meas_start_sr'left);
                i_N_readout_samples <= "000011111";  --32 (one window)
            else
                RAM_rw <= '1';
                RAM_OEb <= '0';
                RAM_ADDR <= RAM_rd_addr;
                meas_peds_ena <= '0';
                i_N_readout_samples <= wave_config_q6.N_readout_samples;
            end if;
        end if;
    end process SRAM_mux;


    ena_logic: process(clk, ped_start_ro, daq_start_ro)
    begin
        if rising_edge(clk) then
            single_bus_ena <= ped_start_ro or daq_start_ro;
        end if;
    end process ena_logic;


    asic_chan_win_mux: process(clk, wave_config_q6.measure_peds, ped_meas_win, daq_asic_mask, trig_q0)
    begin
        if rising_edge(clk) then
            if wave_config_q6.measure_peds = '1' then
                i_trig_bits <= (others=>(others=>'1'));
                asic_mask <= (others=>'1');
                starting_win_samp <= (others=> ped_meas_win & "00000");
                first_dig_win <= ped_meas_win;
                last_dig_win  <= ped_meas_win;
            else
                first_dig_win <= trig_q0.roi_start_addr(10 downto 2);
                last_dig_win  <= trig_q0.roi_stop_addr(10 downto 2);
                asic_mask <= daq_asic_mask;
                for i in 0 to 9 loop
                    starting_win_samp(i) <= (trig_q0.ana_addr(i)(10 downto 0) & "000") - ("00000" & wave_config_q6.ROILookBack & "000");
                    LE_ctime(i) <= (trig_q0.L0_ctime(i)(10 downto 0) & "000") - ("00000" & wave_config_q6.ROILookBack & "000");
                    i_trig_bits(i) <= trig_q0.bits(i); -- used by SingleBusProcessing to make a channel mask
                end loop;
            end if;
        end if;
    end process asic_chan_win_mux;
    ----------------------------------------------------------------------------



    ------------------------------------------------
    --- Process Triggers: Calc ROI, fill queue, mask windows  --  initiated by in port 'localtrg'
    ------------------------------------------------
    trg_proc: process(clk, i_localtrg(i_localtrg'left), queue_full, mask_ack, trig, trg_stg_fsm_ctr)
    begin
        if rising_edge(clk) then
             case trig_staging is
                
                when IDLE =>
                    trg_stg_fsm_ctr <= 0;
                    if i_localtrg(i_localtrg'left) = '1' and queue_full = '0' then  --FIXME: if queue_full=1 or state!=IDLE, then localtrig is ignored
                        trg_proc_busy <= '1';
                        trig_staging <= WAIT_VALID;
                    else
                        trg_proc_busy <= '0';
                        trig_staging <= IDLE;
                    end if;
                
                when WAIT_VALID =>
                    -- tbfifo_rden <= "0000000000";
                    -- if trig.ready = "1111111111" then
                        trig_in_t0 <= trig; -- tb_fifo is 1st-wd fall-through, so trig ready before tbfifo_rden
                        -- tbfifo_rden <= trig.mask;
                        -- tbfifo_rden <= "1111111111"; -- mask taken care of in KLMTrigBitsProc
                        calc_roi_ena <= '1';
                        trig_staging <= PROCESSING_REQ;
                    -- else
                        -- trig_staging <= WAIT_VALID;
                    -- end if;
                
                when PROCESSING_REQ =>
                    -- tbfifo_rden <= "0000000000";
                    calc_roi_ena <= '0';
                    if trg_stg_fsm_ctr < (CALC_ROI_LAG_g + N_ASICS) then
                        trg_stg_fsm_ctr <= trg_stg_fsm_ctr + 1;
                    -- if calc_roi_ena = '1' or calc_roi_busy(1) = '1' or calc_roi_busy(0) = '1' then -- wait for calcROI
                        trig_staging <= PROCESSING_REQ;
                    -- elsif or_calc_roi_busy = '1' then
                    --     trig_staging <= PROCESSING_REQ;
                    else
                        mask_windows <= '1'; -- stop TargetX sampling over ROI
                        trig_queue_wr_ena <= '1'; -- trig_in_t1 ready w/ROI info added. Add to queue.
                        trig_staging <= WAIT_ACK;
                    end if;
                    
                when WAIT_ACK =>
                    trig_queue_wr_ena <= '0';
                    if mask_ack = '1' then -- wait for verification that masking was done
                        mask_windows <= '0';
                        trig_staging <= IDLE;
                    else
                        trig_staging <= WAIT_ACK;
                    end if;

            end case;
        end if;
    end process trg_proc;


    ------------------------------------------------
    --- Queue triggers and initiate readout
    ------------------------------------------------
    trg_queue: process(clk, i_b2tt_runreset, trig_queue_wr_ena, queue_full,
                       queue_empty, hit_bldr_fsm_busy, trig_in_t1)
    begin
        if rising_edge(clk) then
            -- queue_above_thresh <= queue_getting_full or queue_full;
            if i_b2tt_runreset(i_b2tt_runreset'left) = '1' then
                queue_empty <= '1';
                queue_full <= '0';
                start_readout <= '0';
                rd_ptr <= wr_ptr;
            else
                if wr_ptr = (TRIG_QUEUE_DEPTH_g - 1) then
                    wr_ptr_nxt <= 0;
                else
                    wr_ptr_nxt <= wr_ptr + 1;
                end if;
                -- if wr_ptr >= rd_ptr then
                --     if (wr_ptr - rd_ptr) >= TQ_PROG_FULL_THRESH_g then
                --         queue_getting_full <= '1';
                --     else
                --         queue_getting_full <= '0';
                --     end if;
                -- else
                --     if (TRIG_QUEUE_DEPTH_g - (rd_ptr - wr_ptr)) >= TQ_PROG_FULL_THRESH_g then
                --         queue_getting_full <= '1';
                --     else
                --         queue_getting_full <= '0';
                --     end if;
                -- end if;
                if rd_ptr = (TRIG_QUEUE_DEPTH_g - 1) then
                    rd_ptr_nxt <= 0;
                else
                    rd_ptr_nxt <= rd_ptr + 1;
                end if;
                if trig_queue_wr_ena = '1' and queue_full = '0'then
                    trig_queue(wr_ptr) <= trig_in_t1; -- Add trigger to queue
                    if wr_ptr = (TRIG_QUEUE_DEPTH_g - 1) then -- increment write pointer
                        wr_ptr <= 0;
                    else
                        wr_ptr <= wr_ptr + 1;
                    end if;
                    if wr_ptr_nxt = rd_ptr then
                        queue_full <= '1';
                    end if;
                    queue_empty <= '0';
                elsif queue_empty = '0' and hit_bldr_fsm_busy = '0' and start_readout = '0' then
                    start_readout <= '1'; -- initiate readout
                    trig_q0 <= trig_queue(rd_ptr); -- trig_q0 is the one being processed
                    if rd_ptr = (TRIG_QUEUE_DEPTH_g - 1) then -- increment read pointer
                        rd_ptr <= 0;
                    else
                        rd_ptr <= rd_ptr + 1;
                    end if;
                    if rd_ptr_nxt = wr_ptr then
                        queue_empty <= '1';
                    end if; 
                    queue_full <= '0';
                else
                    start_readout <= '0';
                end if;
            end if;
        end if;
    end process trg_queue;


    ------------------------------------------------
    --- Mask / Unmask windows for waveform sampling
    ------------------------------------------------
    mask_unmask_proc: process(clk, mask_windows, unmask_windows, mod_samp_msk_fsm_ctr,
                              trig_in_t1.roi_start_addr, trig_q0.roi_start_addr)
    begin
        if rising_edge(clk) then
            case modify_sampling_mask is
            
                when IDLE =>
                    mod_samp_msk_fsm_ctr <= 0;
                    i_ana_wr_ena_mask <= null_TX_ana_wr_ena_mask;
                    mask_ack <= '0';
                    unmask_ack <= '0';
                    if mask_windows = '1' then -- mask off windows when trigger goes into queue (trig_in_t1)
                        mask_ack <= '1'; -- acknowledge signal to arbitrate collisions
                        i_ana_wr_ena_mask.ena <= trig_in_t1.is_hit;
                        i_ana_wr_ena_mask.mask_bit <= '0';
                        i_ana_wr_ena_mask.win_start <= trig_in_t1.roi_start_addr(10 downto 2);
                        i_ana_wr_ena_mask.n_win <= trig_in_t1.roi_width;
                        modify_sampling_mask <= WAIT_DONE;
                    elsif unmask_windows = '1' then -- unmask windows when current trigger (trig_q0) is done processing
                        unmask_ack <= '1';
                        i_ana_wr_ena_mask.ena <= trig_q0.is_hit;
                        i_ana_wr_ena_mask.mask_bit <= '1';
                        i_ana_wr_ena_mask.win_start <= trig_q0.roi_start_addr(10 downto 2);
                        i_ana_wr_ena_mask.n_win <= trig_q0.roi_width;
                        modify_sampling_mask <= WAIT_DONE;
                    else
                        modify_sampling_mask <= IDLE;
                    end if;
                    
                when WAIT_DONE =>
                    mask_ack <= '0';
                    unmask_ack <= '0';
                    -- if mod_samp_msk_fsm_ctr = (N_READOUT_SAMPLES(7 downto 5) + "010") then
                    if mod_samp_msk_fsm_ctr = 3 then
                        i_ana_wr_ena_mask <= null_TX_ana_wr_ena_mask;
                        modify_sampling_mask <= IDLE;
                    else
                        mod_samp_msk_fsm_ctr <= mod_samp_msk_fsm_ctr + 1;
                        modify_sampling_mask <= WAIT_DONE;
                    end if;
            
            end case;
        end if;
    end process;

   -----------------------------------------------------------------------------
   --- KLM Hit Builder -- initiated when HitQueue not empty and this FSM not busy
   -----------------------------------------------------------------------------
    hit_bldr: process(clk, i_b2tt_runreset, start_readout, trig_q0.mask, trig_q0.bits, trig_q0.L0_ctime,
            rx_features_ena, peak, le_time, LE_ctime, daq_chan, i_full_proc_cnt, i_simp_proc_cnt, i_null_proc_cnt,
            last_hit, unmask_ack, wave_config_q6.use_ftsw_trig, wave_config_q6.simple_pkt_mode,
            proc_queue_quick, i_first_hit, i_last_hit, ro_st_fsm_ctr, ser_busy, ser_run_q2, ser_run_q3)
    begin
        if rising_edge(clk) then
            if i_b2tt_runreset(i_b2tt_runreset'left) = '1' then
                ro_state <= IDLE;
                ser_run_q0 <= '0';
                qt_fifo_evt_rdy <= '0';
                ro_reset <= '1';
                proc_queue_quick <= '0';
                i_full_proc_cnt <= (others=>'0');
                i_simp_proc_cnt <= (others=>'0');
                i_null_proc_cnt <= (others=>'0');
            else

                case ro_state is

                    WHEN IDLE =>
                        ro_reset <= '0';
                        ser_run_q0 <= '0';
                        qt_fifo_evt_rdy <= '0';
                        i_first_hit <= '1';
                        daq_chan_base <= (others=>'0');
                        if start_readout = '1' then -- initiated by trig_queue whenever queue is nonempty and readout is not busy
                            
                            ro_st_fsm_ctr <= 0;
                            ro_reset <= '1';
                            hit_bldr_fsm_busy <= '1';
                            ro_state <= WAIT_RESET;
                        else
                            hit_bldr_fsm_busy <= '0';
                            ro_state <= IDLE;
                        end if;

                    -- FIXME: CHECK IF STATE CAN BE REMOVED
                    When WAIT_RESET => -- soft reset to make sure staging fifos are empty before processing new trigger
                        if ro_st_fsm_ctr < 3 then
                            ro_reset <= '1';
                        else
                            ro_reset <= '0';
                        end if;
                        if ro_st_fsm_ctr < T_WAIT_2C_IF_QUEUE_FULL_g then
                            ro_st_fsm_ctr <= ro_st_fsm_ctr + 1;
                            ro_state <= WAIT_RESET;
                        else
                            ro_st_fsm_ctr <= 0;
                            HitData_i.last_hit <= '0';
                            HitData_i.null_hit <= '1';
                            ro_state <= CHECK_VALID;
                        end if;


                    -- wait until event data is valid
                    WHEN CHECK_VALID =>
                        i_last_hit(0) <= not or_reduce(trig_q0.mask(4 downto 0));
                        i_last_hit(1) <= not or_reduce(trig_q0.mask(9 downto 5));
                        daq_asic_mask <= trig_q0.mask;
                        simp_asic_mask <= trig_q0.mask;
                        if or_reduce(trig_q0.mask) = '1' then
                            HitData_i.null_hit <= '0';
                            -- if queue_above_thresh = '0' and wave_config_q6.simple_pkt_mode = '0' then
                            if proc_queue_quick = '0' and wave_config_q6.simple_pkt_mode = '0' then
                                simple_mode_ena <= '0';
                                daq_start_ro <= '1';
                                simp <= '0';
                                i_full_proc_cnt <= i_full_proc_cnt + '1';
                                ro_state <= WAIT_WAVEFORM_READOUT;
                            else
                                simple_mode_ena <= '1';
                                simp <= '1';
                                i_simp_proc_cnt <= i_simp_proc_cnt + '1';
                                ro_state <= SEND_SIMPLE;
                            end if;
                        else
                            i_null_proc_cnt <= i_null_proc_cnt + '1';
                            ro_state <= SEND_HITS;
                        end if;


                    WHEN WAIT_WAVEFORM_READOUT =>
                        daq_start_ro <= '0';
                        if rx_features_ena(0) = '1' then
                            rx_features_ack <= "01";
                            daq_axis_i <= '0';
                            peak_i <= peak(0);
                            -- le_time_c <= le_time(0)(13 downto 5);
                            -- le_time_f <= le_time(0)(4 downto 0);
                            le_time_i <= LE_ctime(daq_asic(0)) + le_time(0);
                            daq_chan_i <= daq_chan(0);
                            L0_ctime_i <=  trig_q0.L0_ctime(daq_asic(0));
                            trig_bits_i <= trig_q0.bits(daq_asic(0));
                            i_last_hit(0) <= last_hit(0); -- BusA last hit
                            ro_state <= SEND_HITS;
                        elsif rx_features_ena(1) = '1' then
                            rx_features_ack <= "10";
                            daq_axis_i <= '1';
                            peak_i <= peak(1);
                            -- le_time_c <= le_time(1)(13 downto 5);
                            -- le_time_f <= le_time(1)(4 downto 0);
                            le_time_i <= LE_ctime(daq_asic(1) + 5) + le_time(1);
                            L0_ctime_i <= trig_q0.L0_ctime(daq_asic(1) + 5);
                            trig_bits_i <= trig_q0.bits(daq_asic(1) + 5);
                            daq_chan_i <= daq_chan(1);
                            i_last_hit(1) <= last_hit(1); -- BusB last hit
                            ro_state <= SEND_HITS;
                        else
                            ro_state <= WAIT_WAVEFORM_READOUT;
                        end if;


                    WHEN SEND_HITS =>
                        if simple_mode_ena = '1' then
                            i_last_hit(0) <= not or_reduce(simp_asic_mask(4 downto 0));
                            i_last_hit(1) <= not or_reduce(simp_asic_mask(9 downto 5));
                        end if;
                        rx_features_ack <= "00";
                        if (ser_busy or ser_run_q2 or ser_run_q3) = '1' then
                            ro_state <= SEND_HITS;
                        else
                            HitData_i.first_hit <= i_first_hit;
                            -- HitData_i.last_hit <= i_last_hit(1) and i_last_hit(0);
                            ser_run_q0 <= wave_config_q6.use_ftsw_trig; -- initiate transaction
                            ro_state <= CHECK_DONE;
                        end if;


                    WHEN CHECK_DONE  =>
                        ser_run_q0 <= '0';
                        i_first_hit <= '0';
                        if i_last_hit(1) = '1' and i_last_hit(0) = '1' THEN
                            HitData_i.last_hit <= '1';
                            unmask_windows <= '1';
                            -- i_trg_proc_cnt <= i_trg_proc_cnt + '1';
                            ro_state <= STOP;
                        else
                            if simple_mode_ena = '1' then
                                ro_state <= SEND_SIMPLE;
                            else
                                ro_state <= WAIT_WAVEFORM_READOUT;
                            end if;
                        end if;


                    WHEN STOP =>
                        if unmask_ack = '1' then -- VERY IMPORTANT: stay here until sampling mask is removed.
                            qt_fifo_evt_rdy <= wave_config_q6.use_ftsw_trig;
                            unmask_windows <= '0';
                            proc_queue_quick <= not queue_empty;
                            ro_state <= IDLE;
                        else
                            ro_state <= STOP;
                        end if;

                    When SEND_SIMPLE =>
                        if ro_st_fsm_ctr < 5 then
                            daq_axis_i <= '0';
                        else
                            daq_axis_i <= '1';
                        end if;
                        if simp_asic_mask(ro_st_fsm_ctr) = '1' or ro_st_fsm_ctr = 9 then
                            trig_bits_i <= trig_q0.bits(ro_st_fsm_ctr);
                            le_time_i <= LE_ctime(ro_st_fsm_ctr) + nominal_LE_sample_number_g;
                            -- le_time_c <= trig_q0.L0_ctime(ro_st_fsm_ctr)(10 downto 2);
                            -- le_time_f <= trig_q0.L0_ctime(ro_st_fsm_ctr)(1 downto 0) & "000";
                            L0_ctime_i <= trig_q0.L0_ctime(ro_st_fsm_ctr);
                            peak_i <= "000000000000";
                            daq_chan_i <= daq_chan_base + ("000" & trig_q0.bits(ro_st_fsm_ctr)(3 downto 0));
                            simp_asic_mask(ro_st_fsm_ctr) <= '0';
                            ro_state <= SEND_HITS;
                        else
                            ro_state <= SEND_SIMPLE;
                        end if;
                        if ro_st_fsm_ctr = 4 then
                            daq_chan_base <= "0000000";
                        else
                            daq_chan_base <= daq_chan_base + "0001111";
                        end if;
                        ro_st_fsm_ctr <= ro_st_fsm_ctr + 1;

                end case;
            end if;
        end if;

    end process hit_bldr;


    ppln_hit_data: process(clk, daq_axis_i, daq_chan_i, trig_q0.L1_ctime, simp, trig_bits_i,
                           le_time_i, peak_i, HitData_i, ser_run_q0, ser_run_q1)
    begin
        if rising_edge(clk) then
            HitData_i.word1 <= packet_type_g & daq_axis_i & daq_chan_i;
            HitData_i.word2 <= L0_ctime_i;
            -- HitData_i.word2 <= trig_q0.L1_ctime;
            HitData_i.word3 <= trig_bits_i & le_time_i(13 downto 3); -- want word3(11:0) to have same resolution in simple and featExt modes.
            -- HitData_i.word3 <= trig_bits_i & le_time_c & le_time_f(4 downto 3); -- want word3(11:0) to have same resolution in simple and featExt modes.
            HitData_i.word4 <= simp & le_time_i(2 downto 0) & peak_i;
            -- HitData_i.word4 <= simp & le_time_f(2 downto 0) & peak_i;
            -- HitData_i.word4 <= '0' & le_time_f(2 downto 0) & peak_i;
            HitData <= HitData_i;
            ser_run_q1 <= ser_run_q0;
            ser_run_q2 <= ser_run_q1;
            ser_run_q3 <= ser_run_q2;
        end if;
    end process;




---------------------BEGIN MODULES ---------------------------------------------
    CALC_ROI: entity work.CalculateROI
    -- generic map (
    --     FINE_LOOKBACK_g => FINE_LOOKBACK_g
    -- )
    port map (
        clk         => clk,
        ena         => calc_roi_ena,
        lookback    => wave_config_q6.ROILookBack,
        roi_size    => wave_config_q6.N_readout_samples(8 downto 3),
        -- busy        => calc_roi_busy(i),
        -- vec_arr     => L0_ctime_win,
        vec_arr     => trig_in_t0.ana_addr,
        arr_mask    => trig_in_t0.mask,
        is_hit      => trig_in_t1.is_hit,
        first_vec   => trig_in_t1.roi_start_addr,
        last_vec    => trig_in_t1.roi_stop_addr,
        roi_width   => trig_in_t1.roi_width
    );


    busA : entity work.SingleBusProcessing
    generic map (
        N_BITS_AVG_g             => N_BITS_AVG_g,
        USE_PULSE_HEIGHT_HIST    => USE_PULSE_HEIGHT_HIST,
        USE_DBG_WAVE_FIFO        => USE_DBG_WAVE_FIFO
    )
    port map (
        -- main inputs
        clk                => clk,
        rst                => single_bus_reset_q1,
        ped_sub_ena        => wave_config_q6.ped_sub_ena,
        disambig_tb5       => disambig_tb5,
        measure_peds       => wave_config_q6.measure_peds,
        stream_peds        => wave_config_q6.stream_peds,
        ena                => single_bus_ena,
        win_samp_start     => starting_win_samp(4 downto 0),
        trig_bits          => i_trig_bits(4 downto 0),
        asic_mask          => asic_mask(4 downto 0),
        first_dig_win      => first_dig_win,
        last_dig_win       => last_dig_win,

        -- pedestal data
        ped_fetch_asic_no  => i_ped_fetch_asic_no(0),
        ped_fetch_chan     => ped_fetch_chan(0),
        ped_win_samp_start => ped_win_samp_start(0),
        ped_fetch_ena      => ped_fetch_ena(0),
        ped_fetch_ack      => ped_fetch_ack(0),
        ped_fifo_wr_asic   => ped_fifo_asic_sel,
        ped_fifo_wr_chan   => ped_fifo_chan_sel,
        ped_fifo_wr_ena    => ped_fifo_wr_ena(0),
        ped_fifo_din       => ped_fifo_din,

        -- wires to/from TargetX
        BUS_RD_ENA         => BUSA_RD_ENA,
        BUS_RAMP           => BUSA_RAMP,
        BUS_CLR            => BUSA_CLR,
        BUS_DO             => BUSA_DO,
        SR_CLR             => BUSA_SR_CLEAR,
        SR_CLK             => SR_CLOCK(4 downto 0),
        SR_SEL             => BUSA_SR_SEL,
        BUS_RD_WINSEL      => BUSA_WINSEL,
        SAMPLESEL          => BUSA_SAMPLESEL,
        SAMPLESEL_ANY      => SAMPLESEL_ANY(4 downto 0),

        -- wires to HitDataSerializer
        rx_features_ack    => rx_features_ack(0),
        rx_features_ena    => rx_features_ena(0),
        last_hit           => last_hit(0),
        peak               => peak(0),
        le_time            => le_time(0),
        daq_chan           => daq_chan(0),
        daq_asic           => daq_asic(0),

        -- SCROD config registers
        ramp_length        => wave_config_q6.ramp_length,
        -- force_test_pattern => wave_config_q6.force_test_pattern,
        t_samp_addr_settle => wave_config_q6.t_samp_addr_settle,
        t_setup_ss_any     => wave_config_q6.t_setup_ss_any,
        t_strobe_settle    => wave_config_q6.t_strobe_settle,
        t_sr_clk_high      => wave_config_q6.t_sr_clk_high,
        t_sr_clk_low       => wave_config_q6.t_sr_clk_low,
        t_sr_clk_strobe    => wave_config_q6.t_sr_clk_strobe,
        N_readout_samples  => i_N_readout_samples,
        LE_time_thresh     => wave_config_q6.LE_time_thresh,

        -- status registers
        debug_we           => debug_wave_we(0),
        debug_wave         => debug_wave_din(0),
        debug_pfull        => wave_config_q6.debug_wave_pfull(0),
        -- DigStoreProcBusy   => DigStoreProcBusy(0),
        DigNShiftBusy      => DigNShiftBusy(0),
        -- DigBusy            => DigBusy(0),
        ShiftOutWinBusy    => ShiftOutWinBusy(0),
        ShiftOutSampBusy   => ShiftOutSampBusy(0),
        -- FeatExtBusy        => FeatExtBusy(0),
        -- PedFetchQueueBusy  => PedFetchQueueBusy(0),

        -- wires for ped calc
        prime_fifos        => prime_fifos,
        summing_ena        => summing_ena,
        avg_peds_ena       => avg_peds_ena,
        avg_peds_busy      => avg_peds_busy(0),
        wr_peds2sram_ena   => wr_peds2sram_ena(0),
        wr_peds2sram_ack   => wr_peds2sram_ack(0),
        even_ped           => even_sample(0),
        odd_ped            => odd_sample(0),
        sram_asic_addr     => sram_asic_addr(0),
        sram_chan_addr     => sram_chan_addr(0),
        sram_samp_addr     => sram_samp_addr(0),
        -- fe_dbg            => wave_stat_i(0).fe_dbg_a,
        sps_reset          => sps_reset_sr(sps_reset_sr'left),
        SPS_hist_rd_addr   => wave_config_q6.SPS_hist_rd_addr(0),
        SPS_hist_rd_data   => SPS_hist_rd_data(0)
);


    busB : entity work.SingleBusProcessing
    generic map (
        N_BITS_AVG_g             => N_BITS_AVG_g,
        USE_PULSE_HEIGHT_HIST    => USE_PULSE_HEIGHT_HIST,
        USE_DBG_WAVE_FIFO        => USE_DBG_WAVE_FIFO
    )
    port map (
        -- main inputs
        clk                => clk,
        rst                => single_bus_reset_q1,
        ped_sub_ena        => wave_config_q6.ped_sub_ena,
        disambig_tb5       => disambig_tb5,
        measure_peds       => wave_config_q6.measure_peds,
        stream_peds        => wave_config_q6.stream_peds,
        ena                => single_bus_ena,
        win_samp_start     => starting_win_samp(9 downto 5),
        trig_bits          => i_trig_bits(9 downto 5),
        asic_mask          => asic_mask(9 downto 5),
        first_dig_win      => first_dig_win,
        last_dig_win       => last_dig_win,

        -- pedestal data
        ped_fetch_asic_no  => i_ped_fetch_asic_no(1),
        ped_fetch_chan     => ped_fetch_chan(1),
        ped_win_samp_start => ped_win_samp_start(1),
        ped_fetch_ena      => ped_fetch_ena(1),
        ped_fetch_ack      => ped_fetch_ack(1),
        ped_fifo_wr_asic   => ped_fifo_asic_sel,
        ped_fifo_wr_chan   => ped_fifo_chan_sel,
        ped_fifo_wr_ena    => ped_fifo_wr_ena(1),
        ped_fifo_din       => ped_fifo_din,

        -- wires to/from TargetX
        BUS_RD_ENA         => BUSB_RD_ENA,
        BUS_RAMP           => BUSB_RAMP,
        BUS_CLR            => BUSB_CLR,
        BUS_DO             => BUSB_DO,
        SR_CLR             => BUSB_SR_CLEAR,
        SR_CLK             => SR_CLOCK(9 downto 5),
        SR_SEL             => BUSB_SR_SEL,
        BUS_RD_WINSEL      => BUSB_WINSEL,
        SAMPLESEL          => BUSB_SAMPLESEL,
        SAMPLESEL_ANY      => SAMPLESEL_ANY(9 downto 5),

        -- wires to HitDataSerializer
        rx_features_ack    => rx_features_ack(1),
        rx_features_ena    => rx_features_ena(1),
        last_hit           => last_hit(1),
        peak               => peak(1),
        le_time            => le_time(1),
        daq_chan           => daq_chan(1),
        daq_asic           => daq_asic(1),

        -- SCROD config registers
        ramp_length        => wave_config_q6.ramp_length,
        -- force_test_pattern => wave_config_q6.force_test_pattern,
        t_samp_addr_settle => wave_config_q6.t_samp_addr_settle,
        t_setup_ss_any     => wave_config_q6.t_setup_ss_any,
        t_strobe_settle    => wave_config_q6.t_strobe_settle,
        t_sr_clk_high      => wave_config_q6.t_sr_clk_high,
        t_sr_clk_low       => wave_config_q6.t_sr_clk_low,
        t_sr_clk_strobe    => wave_config_q6.t_sr_clk_strobe,
        N_readout_samples  => i_N_readout_samples,
        LE_time_thresh     => wave_config_q6.LE_time_thresh,

        -- status registers
        debug_we           => debug_wave_we(1),
        debug_wave         => debug_wave_din(1),
        debug_pfull        => wave_config_q6.debug_wave_pfull(1),
        -- DigStoreProcBusy   => DigStoreProcBusy(1),
        DigNShiftBusy      => DigNShiftBusy(1),
        -- DigBusy            => DigBusy(1),
        ShiftOutWinBusy    => ShiftOutWinBusy(1),
        ShiftOutSampBusy   => ShiftOutSampBusy(1),
        -- FeatExtBusy        => FeatExtBusy(1),
        -- PedFetchQueueBusy  => PedFetchQueueBusy(1),

        -- wires for ped calc
        prime_fifos        => prime_fifos,
        summing_ena        => summing_ena,
        avg_peds_ena       => avg_peds_ena,
        avg_peds_busy      => avg_peds_busy(1),
        wr_peds2sram_ena   => wr_peds2sram_ena(1),
        wr_peds2sram_ack   => wr_peds2sram_ack(1),
        even_ped           => even_sample(1),
        odd_ped            => odd_sample(1),
        sram_asic_addr     => sram_asic_addr(1),
        sram_chan_addr     => sram_chan_addr(1),
        sram_samp_addr     => sram_samp_addr(1),
        -- fe_dbg            => wave_stat_i(0).fe_dbg_b,
        sps_reset          => sps_reset_sr(sps_reset_sr'left),
        SPS_hist_rd_addr   => wave_config_q6.SPS_hist_rd_addr(1),
        SPS_hist_rd_data   => SPS_hist_rd_data(1)
    );


    ped_fetcher : entity work.PedestalFetcher
    port map (
        clk               => clk,
        rst               => ro_reset,
        ena               => ped_fetch_ena,
        ack               => ped_fetch_ack,
        asic_addr         => i_ped_fetch_asic_no,
        chan_addr         => ped_fetch_chan,
        win_samp_start    => ped_win_samp_start,
        fifo_asic_sel     => ped_fifo_asic_sel, -- fanned out to busA/B, wr_ena controlled
        fifo_chan_sel     => ped_fifo_chan_sel, -- fanned out to busA/B, wr_ena controlled
        ped_fifo_wr_ena   => ped_fifo_wr_ena,   -- slv[1:0]
        ped_fifo_din      => ped_fifo_din,
        N_readout_samples => i_N_readout_samples,
        RAM_do            => RAM_do,
        RAM_ADDR          => RAM_rd_addr
    );


    ped_writer : entity work.PedestalWriter
    port map (
        clk           => clk,
        ena           => wr_peds2sram_ena,
        ack           => wr_peds2sram_ack,
        chan_addr     => sram_chan_addr,
        asic_addr     => sram_asic_addr,
        samp_addr     => sram_samp_addr,
        win_addr      => ped_meas_win,
        even_sample   => even_sample,
        odd_sample    => odd_sample,
        RAM_din       => i_RAM_din,
        RAM_WEb       => i_RAM_WEb,
        RAM_ADDR      => RAM_wr_addr
    );


    ped_measure : entity work.MeasurePeds
    generic map (
        LAST_WINDOW_ADDRESS => LAST_WINDOW_ADDRESS,
        N_BITS_AVG_g => N_BITS_AVG_g
    )
    port map (
        clk                 => clk,
        ena                 => meas_peds_ena,
        busy                => wave_stat_i(0).ped_meas_busy,
        start_ro            => ped_start_ro,
        trig_win            => ped_meas_win,
        prime_fifos         => prime_fifos,
        summing_ena         => summing_ena,
        cur_win             => cur_win,
        either_bus_busy     => or_busy_sr(or_busy_sr'left),
        avg_peds_ena        => avg_peds_ena,
        avg_peds_busy       => avg_peds_busy,
        ped_dbg             => wave_stat_i(0).ped_dbg
        -- bus_mask            => ped_bus_mask
    );


   HitData_Serializer_i : entity work.KLMHitDataSerializer
   port map(
      clk          => clk,
      rst          => i_b2tt_runreset(i_b2tt_runreset'left),
      run          => ser_run_q2,

      -- daq data to be serialized
      first_hit    => HitData.first_hit, -- hit is the first hit in the event
      last_hit     => HitData.last_hit,  -- hit is the last hit in the event
      null_hit     => HitData.null_hit,  -- hit is null
      word1        => HitData.word1,     -- in
      word2        => HitData.word2,     -- in
      word3        => HitData.word3,     -- in
      word4        => HitData.word4,     -- in

      -- nxt        => nxt,
      fifo_empty   => qt_fifo_empty,
      -- fifo_full  => open,
      fifo_dout    => qt_fifo_dout,
      fifo_ren     => qt_fifo_rd_en,
      fifo_err_cnt => qt_fifo_err_cnt,
      busy         => ser_busy
   );


   tristate : for i in 0 to 7 generate
      sda_buff: IOBUF 
         -- generic map(IFD_DELAY_VALUE => "0", DRIVE => 12, SLEW => "SLOW") <-- Default values, uncomment and change if needed
         port map(o => RAM_do(i), io => RAM_IO(i), i => RAM_din(i), t => RAM_rw);
   end generate;


end Behavioral;
